module mem(input logic [7:0]Sbox_data, 
           output logic [7:0]Out) ;


initial begin
		case (Sbox_data)
			8'h0 : Out = 8'h63;
			8'h1 : Out = 8'h7C;
			8'h2 : Out = 8'h77;
			8'h3 : Out = 8'h7B;
			8'h4 : Out = 8'hF2;
			8'h5 : Out = 8'h6B;
			8'h6 : Out = 8'h6F;
			8'h7 : Out = 8'hC5;
			8'h8 : Out = 8'h30;
			8'h9 : Out = 8'h1;
			8'hA : Out = 8'h67;
			8'hB : Out = 8'h2B;
			8'hC : Out = 8'hFE;
			8'hD : Out = 8'hD7;
			8'hE : Out = 8'hAB;
			8'hF : Out = 8'h76;
			8'h10 : Out = 8'hCA;
			8'h11 : Out = 8'h82;
			8'h12 : Out = 8'hC9;
			8'h13 : Out = 8'h7D;
			8'h14 : Out = 8'hFA;
			8'h15 : Out = 8'h59;
			8'h16 : Out = 8'h47;
			8'h17 : Out = 8'hF0;
			8'h18 : Out = 8'hAD;
			8'h19 : Out = 8'hD4;
			8'h1A : Out = 8'hA2;
			8'h1B : Out = 8'hAF;
			8'h1C : Out = 8'h9C;
			8'h1D : Out = 8'hA4;
			8'h1E : Out = 8'h72;
			8'h1F : Out = 8'hC0;
			8'h20 : Out = 8'hB7;
			8'h21 : Out = 8'hFD;
			8'h22 : Out = 8'h93;
			8'h23 : Out = 8'h26;
			8'h24 : Out = 8'h36;
			8'h25 : Out = 8'h3F;
			8'h26 : Out = 8'hF7;
			8'h27 : Out = 8'hCC;
			8'h28 : Out = 8'h34;
			8'h29 : Out = 8'hA5;
			8'h2A : Out = 8'hE5;
			8'h2B : Out = 8'hF1;
			8'h2C : Out = 8'h71;
			8'h2D : Out = 8'hD8;
			8'h2E : Out = 8'h31;
			8'h2F : Out = 8'h15;
			8'h30 : Out = 8'h4;
			8'h31 : Out = 8'hC7;
			8'h32 : Out = 8'h23;
			8'h33 : Out = 8'hC3;
			8'h34 : Out = 8'h18;
			8'h35 : Out = 8'h96;
			8'h36 : Out = 8'h5;
			8'h37 : Out = 8'h9A;
			8'h38 : Out = 8'h7;
			8'h39 : Out = 8'h12;
			8'h3A : Out = 8'h80;
			8'h3B : Out = 8'hE2;
			8'h3C : Out = 8'hEB;
			8'h3D : Out = 8'h27;
			8'h3E : Out = 8'hB2;
			8'h3F : Out = 8'h75;
			8'h40 : Out = 8'h9;
			8'h41 : Out = 8'h83;
			8'h42 : Out = 8'h2C;
			8'h43 : Out = 8'h1A;
			8'h44 : Out = 8'h1B;
			8'h45 : Out = 8'h6E;
			8'h46 : Out = 8'h5A;
			8'h47 : Out = 8'hA0;
			8'h48 : Out = 8'h52;
			8'h49 : Out = 8'h3B;
			8'h4A : Out = 8'hD6;
			8'h4B : Out = 8'hB3;
			8'h4C : Out = 8'h29;
			8'h4D : Out = 8'hE3;
			8'h4E : Out = 8'h2F;
			8'h4F : Out = 8'h84;
			8'h50 : Out = 8'h53;
			8'h51 : Out = 8'hD1;
			8'h52 : Out = 8'h0;
			8'h53 : Out = 8'hED;
			8'h54 : Out = 8'h20;
			8'h55 : Out = 8'hFC;
			8'h56 : Out = 8'hB1;
			8'h57 : Out = 8'h5B;
			8'h58 : Out = 8'h6A;
			8'h59 : Out = 8'hCB;
			8'h5A : Out = 8'hBE;
			8'h5B : Out = 8'h39;
			8'h5C : Out = 8'h4A;
			8'h5D : Out = 8'h4C;
			8'h5E : Out = 8'h58;
			8'h5F : Out = 8'hCF;
			8'h60 : Out = 8'hD0;
			8'h61 : Out = 8'hEF;
			8'h62 : Out = 8'hAA;
			8'h63 : Out = 8'hFB;
			8'h64 : Out = 8'h43;
			8'h65 : Out = 8'h4D;
			8'h66 : Out = 8'h33;
			8'h67 : Out = 8'h85;
			8'h68 : Out = 8'h45;
			8'h69 : Out = 8'hF9;
			8'h6A : Out = 8'h2;
			8'h6B : Out = 8'h7F;
			8'h6C : Out = 8'h50;
			8'h6D : Out = 8'h3C;
			8'h6E : Out = 8'h9F;
			8'h6F : Out = 8'hA8;
			8'h70 : Out = 8'h51;
			8'h71 : Out = 8'hA3;
			8'h72 : Out = 8'h40;
			8'h73 : Out = 8'h8F;
			8'h74 : Out = 8'h92;
			8'h75 : Out = 8'h9D;
			8'h76 : Out = 8'h38;
			8'h77 : Out = 8'hF5;
			8'h78 : Out = 8'hBC;
			8'h79 : Out = 8'hB6;
			8'h7A : Out = 8'hDA;
			8'h7B : Out = 8'h21;
			8'h7C : Out = 8'h10;
			8'h7D : Out = 8'hFF;
			8'h7E : Out = 8'hF3;
			8'h7F : Out = 8'hD2;
			8'h80 : Out = 8'hCD;
			8'h81 : Out = 8'hC;
			8'h82 : Out = 8'h13;
			8'h83 : Out = 8'hEC;
			8'h84 : Out = 8'h5F;
			8'h85 : Out = 8'h97;
			8'h86 : Out = 8'h44;
			8'h87 : Out = 8'h17;
			8'h88 : Out = 8'hC4;
			8'h89 : Out = 8'hA7;
			8'h8A : Out = 8'h7E;
			8'h8B : Out = 8'h3D;
			8'h8C : Out = 8'h64;
			8'h8D : Out = 8'h5D;
			8'h8E : Out = 8'h19;
			8'h8F : Out = 8'h73;
			8'h90 : Out = 8'h60;
			8'h91 : Out = 8'h81;
			8'h92 : Out = 8'h4F;
			8'h93 : Out = 8'hDC;
			8'h94 : Out = 8'h22;
			8'h95 : Out = 8'h2A;
			8'h96 : Out = 8'h90;
			8'h97 : Out = 8'h88;
			8'h98 : Out = 8'h46;
			8'h99 : Out = 8'hEE;
			8'h9A : Out = 8'hB8;
			8'h9B : Out = 8'h14;
			8'h9C : Out = 8'hDE;
			8'h9D : Out = 8'h5E;
			8'h9E : Out = 8'hB;
			8'h9F : Out = 8'hDB;
			8'hA0 : Out = 8'hE0;
			8'hA1 : Out = 8'h32;
			8'hA2 : Out = 8'h3A;
			8'hA3 : Out = 8'hA;
			8'hA4 : Out = 8'h49;
			8'hA5 : Out = 8'h6;
			8'hA6 : Out = 8'h24;
			8'hA7 : Out = 8'h5C;
			8'hA8 : Out = 8'hC2;
			8'hA9 : Out = 8'hD3;
			8'hAA : Out = 8'hAC;
			8'hAB : Out = 8'h62;
			8'hAC : Out = 8'h91;
			8'hAD : Out = 8'h95;
			8'hAE : Out = 8'hE4;
			8'hAF : Out = 8'h79;
			8'hB0 : Out = 8'hE7;
			8'hB1 : Out = 8'hC8;
			8'hB2 : Out = 8'h37;
			8'hB3 : Out = 8'h6D;
			8'hB4 : Out = 8'h8D;
			8'hB5 : Out = 8'hD5;
			8'hB6 : Out = 8'h4E;
			8'hB7 : Out = 8'hA9;
			8'hB8 : Out = 8'h6C;
			8'hB9 : Out = 8'h56;
			8'hBA : Out = 8'hF4;
			8'hBB : Out = 8'hEA;
			8'hBC : Out = 8'h65;
			8'hBD : Out = 8'h7A;
			8'hBE : Out = 8'hAE;
			8'hBF : Out = 8'h8;
			8'hC0 : Out = 8'hBA;
			8'hC1 : Out = 8'h78;
			8'hC2 : Out = 8'h25;
			8'hC3 : Out = 8'h2E;
			8'hC4 : Out = 8'h1C;
			8'hC5 : Out = 8'hA6;
			8'hC6 : Out = 8'hB4;
			8'hC7 : Out = 8'hC6;
			8'hC8 : Out = 8'hE8;
			8'hC9 : Out = 8'hDD;
			8'hCA : Out = 8'h74;
			8'hCB : Out = 8'h1F;
			8'hCC : Out = 8'h4B;
			8'hCD : Out = 8'hBD;
			8'hCE : Out = 8'h8B;
			8'hCF : Out = 8'h8A;
			8'hD0 : Out = 8'h70;
			8'hD1 : Out = 8'h3E;
			8'hD2 : Out = 8'hB5;
			8'hD3 : Out = 8'h66;
			8'hD4 : Out = 8'h48;
			8'hD5 : Out = 8'h3;
			8'hD6 : Out = 8'hF6;
			8'hD7 : Out = 8'hE;
			8'hD8 : Out = 8'h61;
			8'hD9 : Out = 8'h35;
			8'hDA : Out = 8'h57;
			8'hDB : Out = 8'hB9;
			8'hDC : Out = 8'h86;
			8'hDD : Out = 8'hC1;
			8'hDE : Out = 8'h1D;
			8'hDF : Out = 8'h9E;
			8'hE0 : Out = 8'hE1;
			8'hE1 : Out = 8'hF8;
			8'hE2 : Out = 8'h98;
			8'hE3 : Out = 8'h11;
			8'hE4 : Out = 8'h69;
			8'hE5 : Out = 8'hD9;
			8'hE6 : Out = 8'h8E;
			8'hE7 : Out = 8'h94;
			8'hE8 : Out = 8'h9B;
			8'hE9 : Out = 8'h1E;
			8'hEA : Out = 8'h87;
			8'hEB : Out = 8'hE9;
			8'hEC : Out = 8'hCE;
			8'hED : Out = 8'h55;
			8'hEE : Out = 8'h28;
			8'hEF : Out = 8'hDF;
			8'hF0 : Out = 8'h8C;
			8'hF1 : Out = 8'hA1;
			8'hF2 : Out = 8'h89;
			8'hF3 : Out = 8'hD;
			8'hF4 : Out = 8'hBF;
			8'hF5 : Out = 8'hE6;
			8'hF6 : Out = 8'h42;
			8'hF7 : Out = 8'h68;
			8'hF8 : Out = 8'h41;
			8'hF9 : Out = 8'h99;
			8'hFA : Out = 8'h2D;
			8'hFB : Out = 8'hF;
			8'hFC : Out = 8'hB0;
			8'hFD : Out = 8'h54;
			8'hFE : Out = 8'hBB;
			8'hFF : Out = 8'h16;
			default : Out = 8'h0;
		endcase
	end
	
endmodule












